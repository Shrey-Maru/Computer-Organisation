`include "alu.v"

module test;
reg [31:0] ins,a,b;
reg clk, r, i, j;
wire [31:0] out;
wire branch;

ALU a1(ins,a,b,r,i,j,out,branch);

// always #5 clk = ~clk;

initial begin
    clk = 0;
    $dumpfile("test.vcd");
    $dumpvars(0,test);

    //add
    ins = 32'b00000001010010110100100000100000;
    a =   32'b00000000000000000000000000001010;
    b =   32'b00000000000000000000000000000101;
    r=1;
    i=0;
    j=0;
    #10 $display("c = %b",out);
    //or
    ins = 32'b00000001010010110100100000100101;
    a =   32'b00000000000000000000000000001010;
    b =   32'b00000000000000000000000000010001;
    r=1;
    i=0;
    j=1;
    #10 $display("c = %b",out);


    ins = 32'b00100001010010110000000000000100;
    a =   32'b00000000000000000000000000000010;
    b =   32'b00000000000000000000000000000000;
    r=0;
    i=1;
    j=0;
    #10$display("c = %b",out);

    ins = 32'b00010101010010110100100000100100;
    a =   32'b00000000000000000000000000000010;
    b =   32'b00000000000000000000000000000001;
    r=0;
    i=0;
    j=1;
    #10 $display("branch = %b",branch);

    ins = 32'b00010101010010110100100000100100;
    a =   32'b00000000000000000000000000000010;
    b =   32'b00000000000000000000000000000001;
    r=0;
    i=0;
    j=1;
    #10 $display("branch = %b",branch);

    ins = 32'b00010101010010110100100000100100;
    a =   32'b00000000000000000000000000000010;
    b =   32'b00000000000000000000000000000001;
    r=0;
    i=0;
    j=1;
    #10 $display("branch = %b",branch);

    ins = 32'b00010101010010110100100000100100;
    a =   32'b00000000000000000000000000000010;
    b =   32'b00000000000000000000000000000001;
    r=0;
    i=0;
    j=1;
    #10 $display("branch = %b",branch);



    $finish;
end
endmodule